library ieee;
use ieee.std_logic_1164.all;

entity vhdl_top is
  port(a, b : in  std_logic;
       y    : out std_logic);
end entity;

architecture rtl of vhdl_top is
begin
  y <= a and b;
end architecture;
